module Adder(
input [63:0] A, B,
 output [63:0] Out
 );
 
 assign Out= A+B;
 
 
 endmodule